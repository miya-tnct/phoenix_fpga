
module controller (
	clk_clk,
	led0_pio,
	led1_pio,
	led2_pio,
	led3_pio,
	led4_pio,
	reset_reset_n);	

	input		clk_clk;
	output		led0_pio;
	output		led1_pio;
	output		led2_pio;
	output		led3_pio;
	output		led4_pio;
	input		reset_reset_n;
endmodule
