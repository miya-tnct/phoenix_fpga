module pio_source
(
  input wire pio_in,
  output wire pio_out
);

assign pio_out = 1;//pio_in;

endmodule