module phoenix_fpga
(
  input	clk_25mhz
);

endmodule