// controller.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module controller (
		input  wire  clk_clk,       //   clk.clk
		output wire  led0_pio,      //  led0.pio
		output wire  led1_pio,      //  led1.pio
		output wire  led2_pio,      //  led2.pio
		output wire  led3_pio,      //  led3.pio
		output wire  led4_pio,      //  led4.pio
		input  wire  reset_reset_n  // reset.reset_n
	);

	pio_source led0 (
		.pio_in  (),         //  pio_in.pio
		.pio_out (led0_pio)  // pio_out.pio
	);

	pio_source led1 (
		.pio_in  (),         //  pio_in.pio
		.pio_out (led1_pio)  // pio_out.pio
	);

	pio_source led2 (
		.pio_in  (),         //  pio_in.pio
		.pio_out (led2_pio)  // pio_out.pio
	);

	pio_source led3 (
		.pio_in  (),         //  pio_in.pio
		.pio_out (led3_pio)  // pio_out.pio
	);

	pio_source led4 (
		.pio_in  (),         //  pio_in.pio
		.pio_out (led4_pio)  // pio_out.pio
	);

endmodule
