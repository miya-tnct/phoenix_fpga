module phoenix_fpga ();

endmodule