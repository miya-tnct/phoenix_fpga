module phoenix_fpga
(
  input	clk_25mhz,
  output [4:0] leds
);

endmodule