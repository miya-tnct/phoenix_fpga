module pio_source
(
  input wire pio_in,
  output wire pio_out
);

assign pio_out = pio_in;

endmodule