
module controller (
	clk_clk,
	reset_reset_n,
	led0_pio,
	led1_pio,
	led2_pio,
	led3_pio,
	led4_pio);	

	input		clk_clk;
	input		reset_reset_n;
	output		led0_pio;
	output		led1_pio;
	output		led2_pio;
	output		led3_pio;
	output		led4_pio;
endmodule
